// 64QAM DeModulation
module ofdm_demodulation #(
) (
);

endmodulation
