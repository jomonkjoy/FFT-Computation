module fft_controller #(
) (
);

endmodule
