module fft_compute #(
) (
);

endmodule
