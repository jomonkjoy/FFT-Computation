module fft_N_point_core #(
) (
);

endmdoule
