//* magnitude ~= alpha * max(|I|, |Q|) + beta * min(|I|, |Q|) */
module fft_complex_magnitude (
);

endmodule
