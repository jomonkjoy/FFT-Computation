// mux/demux design for 2048 point FFT Core
module fft_mux_2048x1 #(
) (
);

endmodule
