module fft_n_point_core #(
) (
);

endmodule
